** Profile: "SCHEMATIC1-sim_cuad1_param"  [ C:\Cadence\PSD_14.2\tools\cheby_cuad1-schematic1-sim_cuad1_param.sim ] 

** Creating circuit file "cheby_cuad1-schematic1-sim_cuad1_param.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Cadence\PSD_14.2\tools\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 100 0.1 10Meg
.STEP LIN PARAM R3 1k 3k 0.1k 
.PROBE V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC ".\cheby_cuad1-SCHEMATIC1.net" 


.END
