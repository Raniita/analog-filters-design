** Profile: "SCHEMATIC1-sim_cuad2"  [ C:\Cadence\PSD_14.2\tools\cheby_cuad2-schematic1-sim_cuad2.sim ] 

** Creating circuit file "cheby_cuad2-schematic1-sim_cuad2.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Cadence\PSD_14.2\tools\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 100000 0.1 10Meg
.PROBE V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC ".\cheby_cuad2-SCHEMATIC1.net" 


.END
