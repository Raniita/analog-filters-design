** Profile: "SCHEMATIC1-sim_lineal"  [ C:\Cadence\PSD_14.2\tools\cheby_lineal-schematic1-sim_lineal.sim ] 

** Creating circuit file "cheby_lineal-schematic1-sim_lineal.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Cadence\PSD_14.2\tools\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 10000 0.1 1Meg
.PROBE V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC ".\cheby_lineal-SCHEMATIC1.net" 


.END
