** Profile: "SCHEMATIC1-sim_cuad2_param"  [ C:\Cadence\PSD_14.2\tools\cheby_cuad2-schematic1-sim_cuad2_param.sim ] 

** Creating circuit file "cheby_cuad2-schematic1-sim_cuad2_param.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Cadence\PSD_14.2\tools\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 10000 0.1 10Meg
.STEP LIN PARAM R8 8k 11k 0.2k 
.PROBE V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC ".\cheby_cuad2-SCHEMATIC1.net" 


.END
